// megafunction wizard: %ALTTEMP_SENSE%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTTEMP_SENSE 

// ============================================================
// File Name: s5_alttemp_sense.v
// Megafunction Name(s):
// 			ALTTEMP_SENSE
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.1 Build 177 11/07/2012 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module s5_alttemp_sense (
	ce,
	clk,
	clr,
	tsdcaldone,
	tsdcalo)/* synthesis synthesis_clearbox = 1 */;

	input	  ce;
	input	  clk;
	input	  clr;
	output	  tsdcaldone;
	output	[7:0]  tsdcalo;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: CONSTANT: CLK_FREQUENCY STRING "53.125"
// Retrieval info: CONSTANT: CLOCK_DIVIDER_ENABLE STRING "ON"
// Retrieval info: CONSTANT: CLOCK_DIVIDER_VALUE NUMERIC "80"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "alttemp_sense"
// Retrieval info: CONSTANT: NUMBER_OF_SAMPLES NUMERIC "128"
// Retrieval info: CONSTANT: POI_CAL_TEMPERATURE NUMERIC "85"
// Retrieval info: CONSTANT: SIM_TSDCALO NUMERIC "0"
// Retrieval info: CONSTANT: USER_OFFSET_ENABLE STRING "off"
// Retrieval info: CONSTANT: USE_WYS STRING "on"
// Retrieval info: USED_PORT: ce 0 0 0 0 INPUT NODEFVAL "ce"
// Retrieval info: CONNECT: @ce 0 0 0 0 ce 0 0 0 0
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: USED_PORT: clr 0 0 0 0 INPUT NODEFVAL "clr"
// Retrieval info: CONNECT: @clr 0 0 0 0 clr 0 0 0 0
// Retrieval info: USED_PORT: tsdcaldone 0 0 0 0 OUTPUT NODEFVAL "tsdcaldone"
// Retrieval info: CONNECT: tsdcaldone 0 0 0 0 @tsdcaldone 0 0 0 0
// Retrieval info: USED_PORT: tsdcalo 0 0 8 0 OUTPUT NODEFVAL "tsdcalo[7..0]"
// Retrieval info: CONNECT: tsdcalo 0 0 8 0 @tsdcalo 0 0 8 0
// Retrieval info: GEN_FILE: TYPE_NORMAL s5_alttemp_sense.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL s5_alttemp_sense.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL s5_alttemp_sense.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL s5_alttemp_sense_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL s5_alttemp_sense_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL s5_alttemp_sense.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL s5_alttemp_sense.cmp TRUE TRUE
